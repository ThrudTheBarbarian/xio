///////////////////////////////////////////////////////////////////////////////
// Useful stuff shared across modules
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns

//`default_nettype 	none		// Try to catch error early...

`define OP_NONE		2'b00
`define OP_ADD		2'b01
`define OP_DEL		2'b10

